module top (
    
)